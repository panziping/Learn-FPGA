module data_handle(
	



);

	input clk;
	input rst_n;
	
	input [11:0] adc_data;
	input adc_data_valid_go;

	
	
	
	
	output 
	
	
	
	
	


endmodule